version https://git-lfs.github.com/spec/v1
oid sha256:ef166b2737519749064392250a202788f85e7c1f3c7eafb6e4caaa8e53e53c6f
size 744
