version https://git-lfs.github.com/spec/v1
oid sha256:96434d9fdd6da713596d69b26defd18c1b929d74c9de6049d788057d8287844f
size 1050
