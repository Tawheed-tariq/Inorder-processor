version https://git-lfs.github.com/spec/v1
oid sha256:72ea08846c1d6cb35d3b3861a13e0a566facec8a5c4979082f5ba689de40b5ec
size 1197
