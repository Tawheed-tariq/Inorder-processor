version https://git-lfs.github.com/spec/v1
oid sha256:3cd78ddac438af85259c5447948bab78bec7bab4ec884e1574ff1911dca77f3e
size 2326
